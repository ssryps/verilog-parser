`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.11.2019 01:34:23
// Design Name: 
// Module Name: if_id
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`ifdef if_id.v
`else
`define if_id.v

`include "defines.v"

module if_id(
    input wire clk --clock,
    input wire rst --reset,
    input wire[5:0] stall,
	input wire     flush,
    input wire[`InstAddrBus] if_pc --in_signal,
    input wire[`InstBus] if_inst  --in_signal,
    output reg[`InstAddrBus] id_pc --out_signal,
    output reg[`InstBus] id_inst --out_signal
    ); --this.if_id
    
    always @ (posedge clk) begin
        if (rst == `RstEnable) begin
            id_pc <= `ZeroWord;
            id_inst <= `ZeroWord;
        end else if (flush == 1'b1) begin
			id_pc <= `ZeroWord;
			id_inst <= `ZeroWord;					
		end else if(stall[1] == `Stop && stall[2] == `NoStop) begin
			id_pc <= `ZeroWord;
			id_inst <= `ZeroWord;	
	    end else if(stall[1] == `NoStop) begin
		    id_pc <= if_pc;
		    id_inst <= if_inst;
		end
    end
endmodule

`endif